@00000000
08 00 00 06 00 00 00 00 00 00 00 00 00 00 00 00 
31 08 00 00 42 00 00 10 8C 08 02 00 00 00 00 00 
21 08 00 01 21 08 00 01 21 08 00 01 21 08 00 01 
21 08 00 01 21 08 00 01 21 08 00 01 21 08 00 01 
21 08 00 01 21 08 00 01 21 08 00 01 21 08 00 01 
21 08 00 01 21 08 00 01 21 08 00 01 21 08 00 01 
21 08 00 01 08 00 00 08 21 08 00 01 
@00000200
00 00 00 01 00 00 FF FF 
